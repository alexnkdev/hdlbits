module top_module (
  input clk,
  input d,
  output q
);

  wire q1_to_2;
  wire q2_to_3;

  my_dff instance1(
    .clk(clk),
    .d(d),
    .q(q1_to_2)
  );

  my_dff instance2(
    .clk(clk),
    .d(q1_to_2),
    .q(q2_to_3)
  );

  my_dff instance3(
    .clk(clk),
    .d(q2_to_3),
    .q(q)
  );

endmodule
